
timeunit 1ps; //It specifies the time unit that all the delay will take in the simulation.
timeprecision 1ps;// It specifies the resolution in the simulation.

module ReceiveData_TB8x8;

parameter DATA_WIDTH=8;

 // Input Ports
bit clk;
bit reset;
bit RX=1;

// Output Ports
wire LOCKEDST;
wire LOCKEDL;
wire LOCKEDCMD_N_DATA;
wire LOCKEDCMD_PREPARE_RET;
wire LOCKEDN;


 ReceiveData DUT


(
	.clk(clk),
	.reset(reset),
	.RX(RX),
	/* Output */
	.LOCKEDST(LOCKEDST),
	.LOCKEDL(LOCKEDL),
	.LOCKEDCMD_N_DATA(LOCKEDCMD_N_DATA),
	.LOCKEDCMD_PREPARE_RET(LOCKEDCMD_PREPARE_RET),
	.LOCKEDN(LOCKEDN)
);


initial // Clock generator
  begin
    forever #2 clk = !clk;
  end


initial begin // reset generator

	//Cant Pop
	#0 reset = 0;
	#40 reset = 1;
	

	/////INSTRUCTION ONE
	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//3
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//1
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//7
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

/////////////////////////////////////////////////////////


////////////////////////////////// INSTRUCTION TWO
	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//2
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//3
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
//////////////////////////////////////////////////////////

///////////////////////////////INSTRUCTION THREE

	/////DATA
	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//5
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//8
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	////////DATA


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//1
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	

	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//7
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//1
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//3
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	
	//8
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;



	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;


	
	//0
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//4
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	///////////56 VALUES AT THIS POINT

	////////////////////////

	//E
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;

	//F	
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;	
	#40 RX=0;
	#40 RX=0;
	#40 RX=0;
	#40 RX=1;
	#40 RX=0;
	#40 RX=1;
	#40 RX=1;
	#40 RX=1;
	

end



endmodule
