
timeunit 1ps; //It specifies the time unit that all the delay will take in the simulation.
timeprecision 1ps;// It specifies the resolution in the simulation.

module ReceiveData_TB;

parameter DATA_WIDTH=8;

 // Input Ports
bit clk;
bit reset;
bit RX=1;

// Output Ports
wire LOCKEDST;
wire LOCKEDL;
wire LOCKEDCMD_N_DATA;
wire LOCKEDCMD_PREPARE_RET;
wire LOCKEDN;


 ReceiveData DUT


(
	.clk(clk),
	.reset(reset),
	.RX(RX),
	/* Output */
	.LOCKEDST(LOCKEDST),
	.LOCKEDL(LOCKEDL),
	.LOCKEDCMD_N_DATA(LOCKEDCMD_N_DATA),
	.LOCKEDCMD_PREPARE_RET(LOCKEDCMD_PREPARE_RET),
	.LOCKEDN(LOCKEDN)
);


initial // Clock generator
  begin
    forever #2 clk = !clk;
  end


initial begin // reset generator

	//Cant Pop
	#0 reset = 0;
	#80 reset = 1;
	

	/////INSTRUCTION ONE
	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//3
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	
	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//1
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//5
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

/////////////////////////////////////////////////////////


////////////////////////////////// INSTRUCTION TWO
	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;


	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//2
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//3
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
//////////////////////////////////////////////////////////

///////////////////////////////INSTRUCTION THREE

	/////DATA
	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//3
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//2
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	////////DATA
	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//1
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//7
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//1
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;


	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//3
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	//8
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;


	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	
	//0
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//4
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	////////////////////////

	//E
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;

	//F	
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;	
	#80 RX=0;
	#80 RX=0;
	#80 RX=0;
	#80 RX=1;
	#80 RX=0;
	#80 RX=1;
	#80 RX=1;
	#80 RX=1;
	
	
	
end



endmodule
